module song_rom (
    input clk,
    input [8:0] addr,
    output reg [15:0] dout
);

    wire [15:0] memory [511:0];

    always @(posedge clk)
        dout <= memory[addr];

    // Song 0 (Addresses 0-127)
    assign memory[0] = {1'b0, 6'd49, 6'd12, 3'd0};
    assign memory[1] = {1'b1, 6'd12, 9'd0};
    assign memory[2] = {1'b0, 6'd51, 6'd12, 3'd0};
    assign memory[3] = {1'b1, 6'd12, 9'd0};
    assign memory[4] = {1'b0, 6'd52, 6'd12, 3'd0};
    assign memory[5] = {1'b1, 6'd12, 9'd0};
    assign memory[6] = {1'b0, 6'd54, 6'd12, 3'd0};
    assign memory[7] = {1'b1, 6'd12, 9'd0};
    assign memory[8] = {1'b0, 6'd56, 6'd12, 3'd0};
    assign memory[9] = {1'b1, 6'd12, 9'd0};
    assign memory[10] = {1'b0, 6'd57, 6'd12, 3'd0};
    assign memory[11] = {1'b1, 6'd12, 9'd0};
    assign memory[12] = {1'b0, 6'd59, 6'd12, 3'd0};
    assign memory[13] = {1'b1, 6'd12, 9'd0};
    assign memory[14] = {1'b0, 6'd13, 6'd12, 3'd0};
    assign memory[15] = {1'b1, 6'd12, 9'd0};
    assign memory[16] = {1'b0, 6'd15, 6'd12, 3'd0};
    assign memory[17] = {1'b1, 6'd12, 9'd0};
    assign memory[18] = {1'b0, 6'd16, 6'd12, 3'd0};
    assign memory[19] = {1'b1, 6'd12, 9'd0};
    assign memory[20] = {1'b0, 6'd18, 6'd12, 3'd0};
    assign memory[21] = {1'b1, 6'd12, 9'd0};
    assign memory[22] = {1'b0, 6'd20, 6'd12, 3'd0};
    assign memory[23] = {1'b1, 6'd12, 9'd0};
    assign memory[24] = {1'b0, 6'd21, 6'd12, 3'd0};
    assign memory[25] = {1'b1, 6'd12, 9'd0};
    assign memory[26] = {1'b0, 6'd23, 6'd12, 3'd0};
    assign memory[27] = {1'b1, 6'd12, 9'd0};
    assign memory[28] = {1'b0, 6'd37, 6'd0, 3'd0};
    assign memory[29] = {1'b1, 6'd0, 9'd0};
    assign memory[30] = {1'b0, 6'd0, 6'd0, 3'd0};

    assign memory[31] = {1'b0, 6'd28, 6'd6, 3'd0}; // C4
    assign memory[32] = {1'b1, 6'd6, 9'd0};
    assign memory[33] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[34] = {1'b1, 6'd6, 9'd0};
    assign memory[35] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[36] = {1'b1, 6'd6, 9'd0};
    assign memory[37] = {1'b0, 6'd40, 6'd6, 3'd0}; // C5
    assign memory[38] = {1'b1, 6'd6, 9'd0};
    assign memory[39] = {1'b0, 6'd28, 6'd6, 3'd0}; // C4
    assign memory[40] = {1'b1, 6'd6, 9'd0};
    assign memory[41] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[42] = {1'b1, 6'd6, 9'd0};
    assign memory[43] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[44] = {1'b1, 6'd6, 9'd0};
    assign memory[45] = {1'b0, 6'd40, 6'd6, 3'd0}; // C5
    assign memory[46] = {1'b1, 6'd6, 9'd0};
    assign memory[47] = {1'b0, 6'd28, 6'd6, 3'd0}; // C4
    assign memory[48] = {1'b1, 6'd6, 9'd0};
    assign memory[49] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[50] = {1'b1, 6'd6, 9'd0};
    assign memory[51] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[52] = {1'b1, 6'd6, 9'd0};
    assign memory[53] = {1'b0, 6'd40, 6'd6, 3'd0}; // C5
    assign memory[54] = {1'b1, 6'd6, 9'd0};
    assign memory[55] = {1'b0, 6'd28, 6'd6, 3'd0}; // C4
    assign memory[56] = {1'b1, 6'd6, 9'd0};
    assign memory[57] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[58] = {1'b1, 6'd6, 9'd0};
    assign memory[59] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[60] = {1'b1, 6'd6, 9'd0};
    assign memory[61] = {1'b0, 6'd40, 6'd6, 3'd0}; // C5
    assign memory[62] = {1'b1, 6'd6, 9'd0};
    assign memory[63] = {1'b0, 6'd30, 6'd6, 3'd0}; // D4
    assign memory[64] = {1'b1, 6'd6, 9'd0};
    assign memory[65] = {1'b0, 6'd33, 6'd6, 3'd0}; // F4
    assign memory[66] = {1'b1, 6'd6, 9'd0};
    assign memory[67] = {1'b0, 6'd37, 6'd6, 3'd0}; // A4
    assign memory[68] = {1'b1, 6'd6, 9'd0};
    assign memory[69] = {1'b0, 6'd42, 6'd6, 3'd0}; // D5
    assign memory[70] = {1'b1, 6'd6, 9'd0};
    assign memory[71] = {1'b0, 6'd30, 6'd6, 3'd0}; // D4
    assign memory[72] = {1'b1, 6'd6, 9'd0};
    assign memory[73] = {1'b0, 6'd33, 6'd6, 3'd0}; // F4
    assign memory[74] = {1'b1, 6'd6, 9'd0};
    assign memory[75] = {1'b0, 6'd37, 6'd6, 3'd0}; // A4
    assign memory[76] = {1'b1, 6'd6, 9'd0};
    assign memory[77] = {1'b0, 6'd42, 6'd6, 3'd0}; // D5
    assign memory[78] = {1'b1, 6'd6, 9'd0};
    assign memory[79] = {1'b0, 6'd30, 6'd6, 3'd0}; // D4
    assign memory[80] = {1'b1, 6'd6, 9'd0};
    assign memory[81] = {1'b0, 6'd33, 6'd6, 3'd0}; // F4
    assign memory[82] = {1'b1, 6'd6, 9'd0};
    assign memory[83] = {1'b0, 6'd37, 6'd6, 3'd0}; // A4
    assign memory[84] = {1'b1, 6'd6, 9'd0};
    assign memory[85] = {1'b0, 6'd42, 6'd6, 3'd0}; // D5
    assign memory[86] = {1'b1, 6'd6, 9'd0};
    assign memory[87] = {1'b0, 6'd30, 6'd6, 3'd0}; // D4
    assign memory[88] = {1'b1, 6'd6, 9'd0};
    assign memory[89] = {1'b0, 6'd33, 6'd6, 3'd0}; // F4
    assign memory[90] = {1'b1, 6'd6, 9'd0};
    assign memory[91] = {1'b0, 6'd37, 6'd6, 3'd0}; // A4
    assign memory[92] = {1'b1, 6'd6, 9'd0};
    assign memory[93] = {1'b0, 6'd42, 6'd6, 3'd0}; // D5
    assign memory[94] = {1'b1, 6'd6, 9'd0};
    assign memory[95] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[96] = {1'b1, 6'd6, 9'd0};
    assign memory[97] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[98] = {1'b1, 6'd6, 9'd0};
    assign memory[99] = {1'b0, 6'd39, 6'd6, 3'd0}; // B4
    assign memory[100] = {1'b1, 6'd6, 9'd0};
    assign memory[101] = {1'b0, 6'd44, 6'd6, 3'd0}; // E5
    assign memory[102] = {1'b1, 6'd6, 9'd0};
    assign memory[103] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[104] = {1'b1, 6'd6, 9'd0};
    assign memory[105] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[106] = {1'b1, 6'd6, 9'd0};
    assign memory[107] = {1'b0, 6'd39, 6'd6, 3'd0}; // B4
    assign memory[108] = {1'b1, 6'd6, 9'd0};
    assign memory[109] = {1'b0, 6'd44, 6'd6, 3'd0}; // E5
    assign memory[110] = {1'b1, 6'd6, 9'd0};
    assign memory[111] = {1'b0, 6'd32, 6'd6, 3'd0}; // E4
    assign memory[112] = {1'b1, 6'd6, 9'd0};
    assign memory[113] = {1'b0, 6'd35, 6'd6, 3'd0}; // G4
    assign memory[114] = {1'b1, 6'd6, 9'd0};
    assign memory[115] = {1'b0, 6'd39, 6'd6, 3'd0}; // B4
    assign memory[116] = {1'b1, 6'd6, 9'd0};
    assign memory[117] = {1'b0, 6'd44, 6'd6, 3'd0}; // E5
    assign memory[118] = {1'b1, 6'd6, 9'd0};
    assign memory[119] = {1'b0, 6'd28, 6'd24, 3'd0}; // C4 Long
    assign memory[120] = {1'b1, 6'd24, 9'd0};
    assign memory[121] = {1'b0, 6'd0, 6'd0, 3'd0};   // End
    
    // Zero Padding to 127
    assign memory[122] = 16'd0;
    assign memory[123] = 16'd0;
    assign memory[124] = 16'd0;
    assign memory[125] = 16'd0;
    assign memory[126] = 16'd0;
    assign memory[127] = 16'd0;

    // Song 1 (Addresses 128-255)
	
    assign memory[128] = {1'b0, 6'd35, 6'd36, 3'd0};
    assign memory[129] = {1'b0, 6'd39, 6'd36, 3'd0}; 
    assign memory[130] = {1'b0, 6'd42, 6'd36, 3'd0}; 
    assign memory[131] = {1'b1, 6'd36, 9'd0};
    assign memory[132] = {1'b0, 6'd38, 6'd54, 3'd0};
    assign memory[133] = {1'b1, 6'd18, 9'd0};
    assign memory[134] = {1'b0, 6'd37, 6'd18, 3'd0};
    assign memory[135] = {1'b1, 6'd18, 9'd0};
    assign memory[136] = {1'b0, 6'd35, 6'd18, 3'd0};
    assign memory[137] = {1'b1, 6'd18, 9'd0};
    assign memory[138] = {1'b0, 6'd38, 6'd18, 3'd0};
    assign memory[139] = {1'b1, 6'd18, 9'd0};
    assign memory[140] = {1'b0, 6'd37, 6'd18, 3'd0};
    assign memory[141] = {1'b1, 6'd18, 9'd0};
    assign memory[142] = {1'b0, 6'd35, 6'd18, 3'd0};
    assign memory[143] = {1'b1, 6'd18, 9'd0};
    assign memory[144] = {1'b0, 6'd34, 6'd18, 3'd0};
    assign memory[145] = {1'b1, 6'd18, 9'd0};
    assign memory[146] = {1'b0, 6'd37, 6'd18, 3'd0};
    assign memory[147] = {1'b1, 6'd18, 9'd0};
    assign memory[148] = {1'b0, 6'd30, 6'd36, 3'd0};
    assign memory[149] = {1'b1, 6'd36, 9'd0};
    assign memory[150] = {1'b0, 6'd35, 6'd18, 3'd0};
    assign memory[151] = {1'b1, 6'd18, 9'd0};
    assign memory[152] = {1'b0, 6'd30, 6'd18, 3'd0};
    assign memory[153] = {1'b1, 6'd18, 9'd0};
    assign memory[154] = {1'b0, 6'd37, 6'd18, 3'd0};
    assign memory[155] = {1'b1, 6'd18, 9'd0};
    assign memory[156] = {1'b0, 6'd30, 6'd18, 3'd0};
    assign memory[157] = {1'b1, 6'd18, 9'd0};
    assign memory[158] = {1'b0, 6'd38, 6'd18, 3'd0};
    assign memory[159] = {1'b1, 6'd18, 9'd0};
    assign memory[160] = {1'b0, 6'd0, 6'd0, 3'd0};

    assign memory[161] = {1'b0, 6'd32, 6'd8, 3'd0}; // E4
    assign memory[162] = {1'b1, 6'd8, 9'd0};
    assign memory[163] = {1'b0, 6'd35, 6'd8, 3'd0}; // G4
    assign memory[164] = {1'b1, 6'd8, 9'd0};
    assign memory[165] = {1'b0, 6'd37, 6'd8, 3'd0}; // A4
    assign memory[166] = {1'b1, 6'd8, 9'd0};
    assign memory[167] = {1'b0, 6'd39, 6'd8, 3'd0}; // B4
    assign memory[168] = {1'b1, 6'd8, 9'd0};
    assign memory[169] = {1'b0, 6'd42, 6'd8, 3'd0}; // D5
    assign memory[170] = {1'b1, 6'd8, 9'd0};
    assign memory[171] = {1'b0, 6'd44, 6'd8, 3'd0}; // E5
    assign memory[172] = {1'b1, 6'd8, 9'd0};
    assign memory[173] = {1'b0, 6'd47, 6'd8, 3'd0}; // G5
    assign memory[174] = {1'b1, 6'd8, 9'd0};
    assign memory[175] = {1'b0, 6'd49, 6'd8, 3'd0}; // A5
    assign memory[176] = {1'b1, 6'd8, 9'd0};
    assign memory[177] = {1'b0, 6'd51, 6'd8, 3'd0}; // B5
    assign memory[178] = {1'b1, 6'd8, 9'd0};
    assign memory[179] = {1'b0, 6'd54, 6'd8, 3'd0}; // D6
    assign memory[180] = {1'b1, 6'd8, 9'd0};
    assign memory[181] = {1'b0, 6'd56, 6'd8, 3'd0}; // E6
    assign memory[182] = {1'b1, 6'd8, 9'd0};
    // Repeat downward
    assign memory[183] = {1'b0, 6'd54, 6'd8, 3'd0};
    assign memory[184] = {1'b1, 6'd8, 9'd0};
    assign memory[185] = {1'b0, 6'd51, 6'd8, 3'd0};
    assign memory[186] = {1'b1, 6'd8, 9'd0};
    assign memory[187] = {1'b0, 6'd49, 6'd8, 3'd0};
    assign memory[188] = {1'b1, 6'd8, 9'd0};
    assign memory[189] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[190] = {1'b1, 6'd8, 9'd0};
    assign memory[191] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[192] = {1'b1, 6'd8, 9'd0};
    assign memory[193] = {1'b0, 6'd42, 6'd8, 3'd0};
    assign memory[194] = {1'b1, 6'd8, 9'd0};
    assign memory[195] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[196] = {1'b1, 6'd8, 9'd0};
    assign memory[197] = {1'b0, 6'd37, 6'd8, 3'd0};
    assign memory[198] = {1'b1, 6'd8, 9'd0};
    assign memory[199] = {1'b0, 6'd35, 6'd8, 3'd0};
    assign memory[200] = {1'b1, 6'd8, 9'd0};
    assign memory[201] = {1'b0, 6'd32, 6'd8, 3'd0};
    assign memory[202] = {1'b1, 6'd8, 9'd0};
    
    // Simple Chord Stabs to finish (Am -> Em)
    assign memory[203] = {1'b0, 6'd37, 6'd12, 3'd0}; // A4
    assign memory[204] = {1'b0, 6'd40, 6'd12, 3'd0}; // C5
    assign memory[205] = {1'b0, 6'd44, 6'd12, 3'd0}; // E5
    assign memory[206] = {1'b1, 6'd12, 9'd0};
    assign memory[207] = {1'b0, 6'd37, 6'd12, 3'd0};
    assign memory[208] = {1'b0, 6'd40, 6'd12, 3'd0};
    assign memory[209] = {1'b0, 6'd44, 6'd12, 3'd0};
    assign memory[210] = {1'b1, 6'd12, 9'd0};
    assign memory[211] = {1'b0, 6'd32, 6'd24, 3'd0}; // E4
    assign memory[212] = {1'b0, 6'd35, 6'd24, 3'd0}; // G4
    assign memory[213] = {1'b0, 6'd39, 6'd24, 3'd0}; // B4
    assign memory[214] = {1'b1, 6'd24, 9'd0};
    assign memory[215] = {1'b0, 6'd0, 6'd0, 3'd0};   // End

    // Song 2 (Addresses 256-383)

    assign memory[256] = {1'b0, 6'd43, 6'd6, 3'd0};
    assign memory[257] = {1'b1, 6'd6, 9'd0};
    assign memory[258] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[259] = {1'b1, 6'd8, 9'd0};
    assign memory[260] = {1'b0, 6'd0, 6'd34, 3'd0};
    assign memory[261] = {1'b1, 6'd34, 9'd0};
    assign memory[262] = {1'b0, 6'd46, 6'd6, 3'd0};
    assign memory[263] = {1'b1, 6'd6, 9'd0};
    assign memory[264] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[265] = {1'b1, 6'd8, 9'd0};
    assign memory[266] = {1'b0, 6'd0, 6'd34, 3'd0};
    assign memory[267] = {1'b1, 6'd34, 9'd0};
    assign memory[268] = {1'b0, 6'd43, 6'd6, 3'd0};
    assign memory[269] = {1'b1, 6'd6, 9'd0};
    assign memory[270] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[271] = {1'b1, 6'd8, 9'd0};
    assign memory[272] = {1'b0, 6'd0, 6'd10, 3'd0};
    assign memory[273] = {1'b1, 6'd10, 9'd0};
    assign memory[274] = {1'b0, 6'd46, 6'd6, 3'd0};
    assign memory[275] = {1'b1, 6'd6, 9'd0};
    assign memory[276] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[277] = {1'b1, 6'd8, 9'd0};
    assign memory[278] = {1'b0, 6'd0, 6'd10, 3'd0};
    assign memory[279] = {1'b1, 6'd10, 9'd0};
    assign memory[280] = {1'b0, 6'd52, 6'd6, 3'd0};
    assign memory[281] = {1'b1, 6'd6, 9'd0};
    assign memory[282] = {1'b0, 6'd51, 6'd8, 3'd0};
    assign memory[283] = {1'b1, 6'd8, 9'd0};
    assign memory[284] = {1'b0, 6'd0, 6'd10, 3'd0};
    assign memory[285] = {1'b1, 6'd10, 9'd0};
    assign memory[286] = {1'b0, 6'd44, 6'd6, 3'd0};
    assign memory[287] = {1'b1, 6'd6, 9'd0};
    assign memory[288] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[289] = {1'b1, 6'd8, 9'd0};
    assign memory[290] = {1'b0, 6'd0, 6'd10, 3'd0};
    assign memory[291] = {1'b1, 6'd10, 9'd0};
    assign memory[292] = {1'b0, 6'd51, 6'd6, 3'd0};
    assign memory[293] = {1'b1, 6'd6, 9'd0};
    assign memory[294] = {1'b0, 6'd50, 6'd56, 3'd0};
    assign memory[295] = {1'b1, 6'd56, 9'd0};
    assign memory[296] = {1'b0, 6'd49, 6'd8, 3'd0};
    assign memory[297] = {1'b1, 6'd8, 9'd0};
    assign memory[298] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[299] = {1'b1, 6'd8, 9'd0};
    assign memory[300] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[301] = {1'b1, 6'd8, 9'd0};
    assign memory[302] = {1'b0, 6'd42, 6'd8, 3'd0};
    assign memory[303] = {1'b1, 6'd8, 9'd0};
    assign memory[304] = {1'b0, 6'd44, 6'd40, 3'd0};
    assign memory[305] = {1'b1, 6'd40, 9'd0};
    assign memory[306] = {1'b0, 6'd0, 6'd0, 3'd0};

    assign memory[307] = {1'b0, 6'd30, 6'd8, 3'd0}; // D4
    assign memory[308] = {1'b1, 6'd8, 9'd0};
    assign memory[309] = {1'b0, 6'd32, 6'd8, 3'd0}; // E4
    assign memory[310] = {1'b1, 6'd8, 9'd0};
    assign memory[311] = {1'b0, 6'd33, 6'd8, 3'd0}; // F4
    assign memory[312] = {1'b1, 6'd8, 9'd0};
    assign memory[313] = {1'b0, 6'd35, 6'd8, 3'd0}; // G4
    assign memory[314] = {1'b1, 6'd8, 9'd0};
    assign memory[315] = {1'b0, 6'd37, 6'd8, 3'd0}; // A4
    assign memory[316] = {1'b1, 6'd8, 9'd0};
    assign memory[317] = {1'b0, 6'd38, 6'd8, 3'd0}; // Bb4
    assign memory[318] = {1'b1, 6'd8, 9'd0};
    assign memory[319] = {1'b0, 6'd40, 6'd8, 3'd0}; // C5
    assign memory[320] = {1'b1, 6'd8, 9'd0};
    assign memory[321] = {1'b0, 6'd42, 6'd8, 3'd0}; // D5
    assign memory[322] = {1'b1, 6'd8, 9'd0};
    // Down
    assign memory[323] = {1'b0, 6'd40, 6'd8, 3'd0};
    assign memory[324] = {1'b1, 6'd8, 9'd0};
    assign memory[325] = {1'b0, 6'd38, 6'd8, 3'd0};
    assign memory[326] = {1'b1, 6'd8, 9'd0};
    assign memory[327] = {1'b0, 6'd37, 6'd8, 3'd0};
    assign memory[328] = {1'b1, 6'd8, 9'd0};
    assign memory[329] = {1'b0, 6'd35, 6'd8, 3'd0};
    assign memory[330] = {1'b1, 6'd8, 9'd0};
    assign memory[331] = {1'b0, 6'd33, 6'd8, 3'd0};
    assign memory[332] = {1'b1, 6'd8, 9'd0};
    assign memory[333] = {1'b0, 6'd32, 6'd8, 3'd0};
    assign memory[334] = {1'b1, 6'd8, 9'd0};
    assign memory[335] = {1'b0, 6'd30, 6'd16, 3'd0}; // D4
    assign memory[336] = {1'b1, 6'd16, 9'd0};
    
    // Final Chord (Dm)
    assign memory[337] = {1'b0, 6'd30, 6'd24, 3'd0};
    assign memory[338] = {1'b0, 6'd33, 6'd24, 3'd0};
    assign memory[339] = {1'b0, 6'd37, 6'd24, 3'd0};
    assign memory[340] = {1'b1, 6'd24, 9'd0};
    assign memory[341] = {1'b0, 6'd0, 6'd0, 3'd0}; // End

    // Song 3 (Addresses 384-511)
    assign memory[384] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[385] = {1'b1, 6'd8, 9'd0};
    assign memory[386] = {1'b0, 6'd45, 6'd8, 3'd0};
    assign memory[387] = {1'b1, 6'd8, 9'd0};
    assign memory[388] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[389] = {1'b1, 6'd8, 9'd0};
    assign memory[390] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[391] = {1'b1, 6'd8, 9'd0};
    assign memory[392] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[393] = {1'b1, 6'd8, 9'd0};
    assign memory[394] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[395] = {1'b1, 6'd8, 9'd0};
    assign memory[396] = {1'b0, 6'd45, 6'd8, 3'd0};
    assign memory[397] = {1'b1, 6'd8, 9'd0};
    assign memory[398] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[399] = {1'b1, 6'd8, 9'd0};
    assign memory[400] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[401] = {1'b1, 6'd8, 9'd0};
    assign memory[402] = {1'b0, 6'd39, 6'd24, 3'd0};
    assign memory[403] = {1'b1, 6'd24, 9'd0};
    assign memory[404] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[405] = {1'b1, 6'd8, 9'd0};
    assign memory[406] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[407] = {1'b1, 6'd8, 9'd0};
    assign memory[408] = {1'b0, 6'd38, 6'd8, 3'd0};
    assign memory[409] = {1'b1, 6'd8, 9'd0};
    assign memory[410] = {1'b0, 6'd45, 6'd8, 3'd0};
    assign memory[411] = {1'b1, 6'd8, 9'd0};
    assign memory[412] = {1'b0, 6'd44, 6'd40, 3'd0};
    assign memory[413] = {1'b1, 6'd40, 9'd0};
    assign memory[414] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[415] = {1'b1, 6'd8, 9'd0};
    assign memory[416] = {1'b0, 6'd45, 6'd8, 3'd0};
    assign memory[417] = {1'b1, 6'd8, 9'd0};
    assign memory[418] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[419] = {1'b1, 6'd8, 9'd0};
    assign memory[420] = {1'b0, 6'd44, 6'd24, 3'd0};
    assign memory[421] = {1'b1, 6'd24, 9'd0};
    assign memory[422] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[423] = {1'b1, 6'd8, 9'd0};
    assign memory[424] = {1'b0, 6'd38, 6'd8, 3'd0};
    assign memory[425] = {1'b1, 6'd8, 9'd0};
    assign memory[426] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[427] = {1'b1, 6'd8, 9'd0};
    assign memory[428] = {1'b0, 6'd44, 6'd24, 3'd0};
    assign memory[429] = {1'b1, 6'd24, 9'd0};
    assign memory[430] = {1'b0, 6'd39, 6'd24, 3'd0};
    assign memory[431] = {1'b1, 6'd24, 9'd0};
    assign memory[432] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[433] = {1'b1, 6'd8, 9'd0};
    assign memory[434] = {1'b0, 6'd38, 6'd8, 3'd0};
    assign memory[435] = {1'b1, 6'd8, 9'd0};
    assign memory[436] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[437] = {1'b1, 6'd8, 9'd0};
    assign memory[438] = {1'b0, 6'd44, 6'd8, 3'd0};
    assign memory[439] = {1'b1, 6'd8, 9'd0};
    assign memory[440] = {1'b0, 6'd39, 6'd48, 3'd0};
    assign memory[441] = {1'b1, 6'd48, 9'd0};
    assign memory[442] = {1'b0, 6'd39, 6'd8, 3'd0};
    assign memory[443] = {1'b1, 6'd8, 9'd0};
    assign memory[444] = {1'b0, 6'd47, 6'd8, 3'd0};
    assign memory[445] = {1'b1, 6'd8, 9'd0};
    assign memory[446] = {1'b0, 6'd0, 6'd0, 3'd0};

    assign memory[447] = {1'b0, 6'd39, 6'd12, 3'd0}; // B4
    assign memory[448] = {1'b1, 6'd12, 9'd0};
    assign memory[449] = {1'b0, 6'd42, 6'd12, 3'd0}; // D5
    assign memory[450] = {1'b1, 6'd12, 9'd0};
    assign memory[451] = {1'b0, 6'd46, 6'd12, 3'd0}; // F#5
    assign memory[452] = {1'b1, 6'd12, 9'd0};
    assign memory[453] = {1'b0, 6'd51, 6'd12, 3'd0}; // B5
    assign memory[454] = {1'b1, 6'd12, 9'd0};
    assign memory[455] = {1'b0, 6'd46, 6'd12, 3'd0}; // F#5
    assign memory[456] = {1'b1, 6'd12, 9'd0};
    assign memory[457] = {1'b0, 6'd42, 6'd12, 3'd0}; // D5
    assign memory[458] = {1'b1, 6'd12, 9'd0};
    assign memory[459] = {1'b0, 6'd39, 6'd24, 3'd0}; // B4 (End on root)
    assign memory[460] = {1'b1, 6'd24, 9'd0};
    assign memory[461] = {1'b0, 6'd0, 6'd0, 3'd0};   // End


endmodule
